// Code your design here
`include "Top.sv"
`include "RegFile.sv"
`include "ProgCtr.sv"
`include "JLUT.sv"
`include "InstROM.sv"
`include "DMem.sv"
`include "Ctrl.sv"
`include "ALU.sv"

